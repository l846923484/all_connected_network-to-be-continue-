// Copyright (C) 1991-2009 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// *****************************************************************************
// This file contains a Verilog test bench template that is freely editable to  
// suit user's needs .Comments are provided in each section to help the user    
// fill out necessary details.                                                  
// *****************************************************************************
// Generated on "04/12/2019 21:33:56"
                                                                                
// Verilog Test Bench template for design : ctrl_1
// 
// Simulation tool : ModelSim (Verilog)
// 

`timescale 1 ps/ 1 ps
module tb_ctrl_1();
// constants                                           
// general purpose registers
reg clk;
reg reset;
reg [15:0] input_data1,input_data2,input_data3,input_data4,
           input_data5,input_data6,input_data7,input_data8,
           input_data9,input_data10,input_data11,input_data12,
           input_data13,input_data14,input_data15,input_data16;
// wires                                               
wire complete1;
wire complete2;
wire [15:0] q1;
wire wren1;

// assign statements (if any)                          
ctrl_1 i1 (
// port map - connection between master ports and signals/registers   
   
	.clk(clk),
	.reset(reset),
	.wren1(wren1),
	.input_data1(input_data1),.input_data2(input_data2),.input_data3(input_data3),.input_data4(input_data4),
   .input_data5(input_data5),.input_data6(input_data6),.input_data7(input_data7),.input_data8(input_data8),
   .input_data9(input_data9),.input_data10(input_data10),.input_data11(input_data11),.input_data12(input_data12),
   .input_data13(input_data13),.input_data14(input_data14),.input_data15(input_data15),.input_data16(input_data16),
	.q1(q1),  
	.complete1(complete1),
	.complete2(complete2)
	
);
initial                                                
begin                                                  
// code that executes only once                        
// insert code here --> begin   
       reset=1'b1;
       input_data1=16'b0000001000000000;  
       input_data2=16'b0000001000000000;  
       input_data3=16'b0000001000000000;  
       input_data4=16'b0000001000000000;  
       input_data5=16'b0000001000000000;  
       input_data6=16'b0000001000000000;  
       input_data7=16'b0000001000000000;  
       input_data8=16'b0000001000000000;  
       input_data9=16'b0000001000000000;  
       input_data10=16'b0000001000000000;  
       input_data11=16'b0000001000000000;  
       input_data12=16'b0000001000000000;  
       input_data13=16'b0000000000000000;  
       input_data14=16'b0000000000000000;  
       input_data15=16'b0000000000000000;  
       input_data16=16'b0000000000000000;     
       #5
       reset=1'b0;                                                      
// --> end                                             
//$display("Running testbench");                       
end     
                                               
initial                     
begin                                           
            clk=1'b0;
            forever #10 clk=~clk;                                                                                  
end                                                    
endmodule

